module And(input a,b output y);
  assign y =a & b;
endmodule
